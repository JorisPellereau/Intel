JorisPC@JORISP.5124:1561451602