JorisPC@JORISP.13860:1561104311