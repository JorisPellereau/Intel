
module NIOS_II_debug (
	clk_clk,
	pio_uart_data_external_connection_export,
	reset_reset_n);	

	input		clk_clk;
	input	[7:0]	pio_uart_data_external_connection_export;
	input		reset_reset_n;
endmodule
